library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity zadatak is
    port (
        A, B: in  STD_LOGIC_VECTOR(1 downto 0);
        C   : out STD_LOGIC_VECTOR(3 downto 0)
    );
end zadatak;

architecture Behavioral of zadatak is
begin
    --------------------------------------------------------------------
    -- C0 = A0 B0
    --------------------------------------------------------------------
    C(0) <= A(0) and B(0);
    --------------------------------------------------------------------
    -- C1 = A1 B0 ⊕ A0 B1
    --------------------------------------------------------------------
    C(1) <= (A(1) and B(0)) xor (A(0) and B(1));
    --------------------------------------------------------------------
    -- C2 = (A1 B1) (A0 nand B0)
    --------------------------------------------------------------------
    C(2) <= (A(1) and B(1)) and (A(0) nand B(0));
    --------------------------------------------------------------------
    -- C3 = A1 A0 B1 B0
    --------------------------------------------------------------------
    C(3) <= A(1) and A(0) and B(1) and B(0);

end Behavioral;