library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity zadatak_4 is
    generic (
        T : time := 1 ns   -- globalni delay parametar
    );
    port (
        A : in  STD_LOGIC;
        B : in  STD_LOGIC;
        C : in  STD_LOGIC;
        D : in  STD_LOGIC;
        Y : out STD_LOGIC
    );
end zadatak_4;

architecture Behavioral of zadatak_4 is
    -- interni signali
    signal B_inv, I1 : STD_LOGIC;
    signal I2, I3, I4 : STD_LOGIC;
begin
    --------------------------------------------------------------------
    -- B_inv = inv B, I1 = inv D
    --------------------------------------------------------------------
    B_inv <= (not B) after T;
    I1    <= (not D) after T;
    --------------------------------------------------------------------
    -- I2 = A B_inv
    --------------------------------------------------------------------
    I2 <= (A and B_inv) after T;
    --------------------------------------------------------------------
    -- I3 = C D
    --------------------------------------------------------------------
    I3 <= (C and D) after T;
    --------------------------------------------------------------------
    -- I4 = A and C and I1   (A C \bar{D})
    --------------------------------------------------------------------
    I4 <= (A and C and I1) after T;
    --------------------------------------------------------------------
    -- Y = I2 + I3 + I4
    --------------------------------------------------------------------
    Y <= (I2 or I3 or I4) after T;

end Behavioral;
